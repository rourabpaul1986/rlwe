ffew
