This component is required for polynomial divider. In current version poly div is part of polynomial divider
