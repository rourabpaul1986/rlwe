Yet to be designed
