yet to be designed
